
module zi_0in_rtld_ctrl_ctrl; 


endmodule 

