module clock_counter(clk,reset_n,out_counterDIV1M);

input clk,reset_n;
output [15:0] out_counterDIV1M;


assign out_counterDIV1M=0;



endmodule
